`include "base_test.sv"
`include "benchmark_test.sv"